 module saida_serial_fd (
    input        clock        ,
    input        reset        ,
    input        proximo      , // Para mandar pegar o proximo digito 
    input        conta        ,
    input        carrega      ,
    input        desloca      ,
    input  [6:0] dados_ascii  ,
    output       saida_serial ,
    output       fim
);
    // fios internos 


    // componentes
  
    
    // Saida serial do transmissor
    assign saida_serial = ;
  
endmodule
